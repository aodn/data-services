netcdf imos_missing_data {
dimensions:
	time = 10 ;
variables:
	double time(time) ;
		time:standard_name = "" ;
		time:valid_min = "" ;
		time:valid_max = "" ;
		time:calendar = "" ;

// global attributes:
		:project = "" ;
		:conventions = "" ;
		:date_created = "" ;
		:geospatial_lat_min = 0L ;
		:geospatial_lat_max = 100L ;
		:naming_authority = "" ;
		:geospatial_lon_min = 0L ;
		:geospatial_lon_max = 100L ;
		:time_coverage_start = 0L ;
		:time_coverage_end = 100L ;
		:data_centre = "" ;
		:author = 123L ;
		:citation = 123L ;
		:long_name = 123L ;
		:acknowledgement = "" ;
		:distribution_statement = "" ;
		:valid_min = 0L ;
		:valid_max = 0L ;
data:

 time = _, _, _, _, _, _, _, _, _, _ ;
}

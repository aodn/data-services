netcdf srs_good_data {
dimensions:
	time = 1 ;
	lat = 11 ;
	lon = 26 ;
variables:
	byte dt_analysis(time, lat, lon) ;
		dt_analysis:_FillValue = -128b ;
		dt_analysis:long_name = "deviation from last SST analysis" ;
		dt_analysis:units = "kelvin" ;
		dt_analysis:coordinates = "time lat lon" ;
		dt_analysis:comment = "The difference between this SST and the previous day\'s SST" ;
		dt_analysis:source = "NCDC-L4LRblend-GLOB-AVHRR_OI" ;
		dt_analysis:add_offset = -1.3220397233963 ;
		dt_analysis:scale_factor = 0.0304610503049707 ;
		dt_analysis:valid_min = -127b ;
		dt_analysis:valid_max = 127b ;
	short l2p_flags(time, lat, lon) ;
		l2p_flags:_FillValue = -32768s ;
		l2p_flags:long_name = "L2P flags" ;
		l2p_flags:valid_min = 0s ;
		l2p_flags:valid_max = 32767s ;
		l2p_flags:coordinates = "time lat lon" ;
		l2p_flags:comment = "These flags are important to properly use the data.  Data not flagged as microwave are sourced from an infrared sensor. The lake and river flags are currently not set, but defined in GDS2.0r4. The aerosol flag indicates high aerosol concentration. The analysis flag indicates high difference from analysis temperatures (differences greater than Analysis Limit). The lowwind flag indicates regions of low wind speed (typically less than the low Wind Limit) per NWP model. The highwind flag indicates regions of high wind speed (typically greater than the high Wind Limit) per NWP model. See wind limits in the comment field for the actual values. The edge flag indicates pixel sizes that are larger than Pixel Spread times the size of the pixel in the center of the field of view in either lat or lon direction. The terminator flag indicates that the sun is near the horizon. The reflector flag indicates that the satellite would receive direct reflected sunlight if the earth was a perfect mirror. The swath flag is used in gridded files to indicate if the pixel could have been seen by the satellite. delta_dn indicates that the day.night sst algorithm was different from the standard algorithm. Other flags may be populated and are for internal use and the definitions may change, so should not be relied on. Flags greater than 64 only apply to non-land pixels" ;
		l2p_flags:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s ;
		l2p_flags:flag_meanings = "microwave land ice lake river reserved aerosol analysis lowwind highwind edge terminator reflector swath delta_dn" ;
	float lat(lat) ;
		lat:_FillValue = 9.96921e+36f ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:axis = "Y" ;
		lat:comment = "Latitudes for locating data" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:_FillValue = 9.96921e+36f ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 360.f ;
		lon:axis = "X" ;
		lon:comment = "Longitudes for locating data" ;
		lon:standard_name = "longitude" ;
	byte quality_level(time, lat, lon) ;
		quality_level:_FillValue = -128b ;
		quality_level:long_name = "quality level of SST pixel" ;
		quality_level:valid_min = 0b ;
		quality_level:valid_max = 5b ;
		quality_level:coordinates = "time lat lon" ;
		quality_level:comment = "These are the overall quality indicators and are used for all GHRSST SSTs. In this case they are a function of distance to cloud, satellite zenith angle, and day/night" ;
		quality_level:flag_meanings = "no_data bad_data worst_quality low_quality acceptable_quality best_quality" ;
		quality_level:flag_values = 0b, 1b, 2b, 3b, 4b, 5b ;
	byte satellite_zenith_angle(time, lat, lon) ;
		satellite_zenith_angle:_FillValue = -128b ;
		satellite_zenith_angle:long_name = "satellite zenith angle" ;
		satellite_zenith_angle:units = "angular_degree" ;
		satellite_zenith_angle:coordinates = "time lat lon" ;
		satellite_zenith_angle:comment = "The satellite zenith angle at the time of the SST observations" ;
		satellite_zenith_angle:add_offset = 35.145679473877 ;
		satellite_zenith_angle:scale_factor = 0.270908491413584 ;
		satellite_zenith_angle:valid_min = -127b ;
		satellite_zenith_angle:valid_max = 127b ;
	byte sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:_FillValue = -128b ;
		sea_ice_fraction:long_name = "sea ice fraction" ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:coordinates = "time lat lon" ;
		sea_ice_fraction:comment = "Fractional sea ice cover (Unitless). For spatial resolution refer to the source." ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:source = "SSMI-NCEP-Analysis-ICE-1deg" ;
		sea_ice_fraction:add_offset = 0.388769209384918 ;
		sea_ice_fraction:scale_factor = 0.00298716004186939 ;
		sea_ice_fraction:valid_min = -127b ;
		sea_ice_fraction:valid_max = 127b ;
	byte sea_ice_fraction_dtime_from_sst(time, lat, lon) ;
		sea_ice_fraction_dtime_from_sst:_FillValue = -128b ;
		sea_ice_fraction_dtime_from_sst:long_name = "time difference of sea ice fraction measurement from sst measurement" ;
		sea_ice_fraction_dtime_from_sst:units = "hour" ;
		sea_ice_fraction_dtime_from_sst:coordinates = "time lat lon" ;
		sea_ice_fraction_dtime_from_sst:comment = "The time difference in hours is estimated from the SST and sea ice data sets" ;
		sea_ice_fraction_dtime_from_sst:source = "SSMI-NCEP-Analysis-ICE-1deg" ;
		sea_ice_fraction_dtime_from_sst:add_offset = 20.3899959661067 ;
		sea_ice_fraction_dtime_from_sst:scale_factor = 0.0138194096300442 ;
		sea_ice_fraction_dtime_from_sst:valid_min = -127b ;
		sea_ice_fraction_dtime_from_sst:valid_max = 127b ;
	short sea_surface_temperature(time, lat, lon) ;
		sea_surface_temperature:_FillValue = -32768s ;
		sea_surface_temperature:long_name = "sea surface skin temperature" ;
		sea_surface_temperature:units = "kelvin" ;
		sea_surface_temperature:coordinates = "time lat lon" ;
		sea_surface_temperature:standard_name = "sea_surface_skin_temperature" ;
		sea_surface_temperature:add_offset = 281.99284362793 ;
		sea_surface_temperature:scale_factor = 0.00999999977648258 ;
		sea_surface_temperature:valid_min = -32767s ;
		sea_surface_temperature:valid_max = 32767s ;
		sea_surface_temperature:comment = "The skin temperature of the ocean at a depth of approximately 10um" ;
	short sea_surface_temperature_day_night(time, lat, lon) ;
		sea_surface_temperature_day_night:_FillValue = -32768s ;
		sea_surface_temperature_day_night:units = "kelvin" ;
		sea_surface_temperature_day_night:coordinates = "time lat lon" ;
		sea_surface_temperature_day_night:add_offset = 281.9990234375 ;
		sea_surface_temperature_day_night:scale_factor = 0.00999999977648258 ;
		sea_surface_temperature_day_night:valid_min = -32767s ;
		sea_surface_temperature_day_night:valid_max = 32767s ;
		sea_surface_temperature_day_night:long_name = "sea surface skin temperature" ;
		sea_surface_temperature_day_night:comment = "The skin temperature of the ocean at a depth of approximately 10um based on a unified day / night model - EXPERIMENTAL" ;
		sea_surface_temperature_day_night:standard_name = "sea_surface_skin_temperature" ;
	byte sses_bias(time, lat, lon) ;
		sses_bias:_FillValue = -128b ;
		sses_bias:long_name = "SSES bias estimate" ;
		sses_bias:units = "kelvin" ;
		sses_bias:coordinates = "time lat lon" ;
		sses_bias:add_offset = -0.614610850811005 ;
		sses_bias:scale_factor = 0.0138956515685372 ;
		sses_bias:valid_min = -127b ;
		sses_bias:valid_max = 127b ;
		sses_bias:comment = "Bias estimate derived from L2P bias per https://www.ghrsst.org/ghrsst/tags-and-wgs/stval-wg/sses-description-of-schemes/" ;
	byte sses_count(time, lat, lon) ;
		sses_count:_FillValue = -128b ;
		sses_count:long_name = "SSES count" ;
		sses_count:units = "count" ;
		sses_count:coordinates = "time lat lon" ;
		sses_count:comment = "Weighted representative number of swath pixels. EXPERIMENTAL_FIELD" ;
		sses_count:add_offset = 3.01456040143967 ;
		sses_count:scale_factor = 0.015627750294953 ;
		sses_count:valid_min = -127b ;
		sses_count:valid_max = 127b ;
	byte sses_standard_deviation(time, lat, lon) ;
		sses_standard_deviation:_FillValue = -128b ;
		sses_standard_deviation:long_name = "SSES standard deviation estimate" ;
		sses_standard_deviation:units = "kelvin" ;
		sses_standard_deviation:coordinates = "time lat lon" ;
		sses_standard_deviation:add_offset = 1.04265016317368 ;
		sses_standard_deviation:scale_factor = 0.00587929331738016 ;
		sses_standard_deviation:valid_min = -127b ;
		sses_standard_deviation:valid_max = 127b ;
		sses_standard_deviation:comment = "Standard deviation estimate derived from L2P standard deviation per https://www.ghrsst.org/ghrsst/tags-and-wgs/stval-wg/sses-description-of-schemes/" ;
	int sst_dtime(time, lat, lon) ;
		sst_dtime:_FillValue = -2147483647 ;
		sst_dtime:long_name = "time difference from reference time" ;
		sst_dtime:units = "second" ;
		sst_dtime:coordinates = "time lat lon" ;
		sst_dtime:comment = "time plus sst_dtime gives seconds after 00:00:00 UTC January 1, 1981" ;
		sst_dtime:add_offset = 18173.2557021081 ;
		sst_dtime:scale_factor = 2.93129655703861e-06 ;
		sst_dtime:valid_min = -2147483645 ;
		sst_dtime:valid_max = 2147483645 ;
	int time(time) ;
		time:_FillValue = -2147483647 ;
		time:long_name = "reference time of sst file" ;
		time:units = "seconds since 1981-01-01 00:00:00" ;
		time:axis = "T" ;
		time:comment = "A typical reference time for data" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
	byte wind_speed(time, lat, lon) ;
		wind_speed:_FillValue = -128b ;
		wind_speed:long_name = "wind speed" ;
		wind_speed:units = "m s-1" ;
		wind_speed:coordinates = "time lat lon" ;
		wind_speed:comment = "Typically represent surface winds (10 meters above the sea surface)" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:source = "ECMWF_interim_reanalysis" ;
		wind_speed:height = "10m" ;
		wind_speed:add_offset = 11.5929851531982 ;
		wind_speed:scale_factor = 0.0841179195600065 ;
		wind_speed:valid_min = -127b ;
		wind_speed:valid_max = 127b ;
	byte wind_speed_dtime_from_sst(time, lat, lon) ;
		wind_speed_dtime_from_sst:_FillValue = -128b ;
		wind_speed_dtime_from_sst:long_name = "time difference of wind speed measurement from sst measurement" ;
		wind_speed_dtime_from_sst:units = "hour" ;
		wind_speed_dtime_from_sst:coordinates = "time lat lon" ;
		wind_speed_dtime_from_sst:comment = "The hours between the wind speed measurement and the SST observation" ;
		wind_speed_dtime_from_sst:source = "ECMWF_interim_reanalysis" ;
		wind_speed_dtime_from_sst:add_offset = 0.273298216983676 ;
		wind_speed_dtime_from_sst:scale_factor = 0.0173675635085982 ;
		wind_speed_dtime_from_sst:valid_min = -127b ;
		wind_speed_dtime_from_sst:valid_max = 127b ;

// global attributes:
		:title = "IMOS L3S Daytime gridded multiple-sensor multiple-swath Australian region HRPT AVHRR skin SST" ;
		:summary = "Skin SST retrievals produced from stitching together High Resolution Picture Transmission direct broadcast data from a NOAA polar-orbiting satellite received at Australian receiving stations." ;
		:institution = "ABOM" ;
		:license = "GHRSST protocol describes data use as free and open" ;
		:id = "AVHRR_D-ABOM-L3S-v02.0" ;
		:naming_authority = "org.ghrsst" ;
		:uuid = "d77fe51d-2fe6-4ad8-a3b4-16b6ea641247" ;
		:gds_version_id = "2.0r4" ;
		:netcdf_version_id = "4.2.1.1" ;
		:date_created = "20141010T075620Z" ;
		:file_quality_level = 3 ;
		:spatial_resolution = "0.02 deg" ;
		:start_time = "19920326T063758Z" ;
		:time_coverage_start = "19920326T063758Z" ;
		:stop_time = "19920326T100748Z" ;
		:time_coverage_end = "19920326T100748Z" ;
		:northernmost_latitude = 19.99f ;
		:southernmost_latitude = -69.99f ;
		:easternmost_longitude = -170.01f ;
		:westernmost_longitude = 70.01f ;
		:source = "wind_source=ECMWF_interim_reanalysis,analysis_source=NCDC-L4LRblend-GLOB-AVHRR_OI,adi_source=unknown,ice_source=SSMI-NCEP-Analysis-ICE-1deg,l3_source=AVHRR11_D-ABOM-L3C-v02.0" ;
		:platform = "NOAA-11" ;
		:sensor = "AVHRR" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:Metadata_Link = "TBA" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = 0.02f ;
		:geospatial_lon_resolution = 0.02f ;
		:creator_name = "Australian Bureau of Meteorology" ;
		:creator_email = "ghrsst@bom.gov.au" ;
		:project = "Group for High Resolution Sea Surface Temperature" ;
		:publisher_name = "The GHRSST Project Office" ;
		:publisher_email = "ghrsst-po@nceo.ac.uk" ;
		:publisher_url = "http://www.ghrsst.org" ;
		:processing_level = "L3S" ;
		:cdm_data_type = "grid" ;
		:history = "Tue Oct 18 16:40:51 2016: ncks -d lat,30,40 -d lon,25,50 data/srs_new_data.nc -O srs_good_data.nc\nplatform_counts=NOAA-11=1,quality_counts=archive=1,platform=NOAA-11,quality_source=archive,ice_source=SSMI-NCEP-Analysis-ICE-1deg,adi_source=unknown,wind_source=ECMWF_interim_reanalysis,analysis_source=NCDC-L4LRblend-GLOB-AVHRR_OI,source_file=19920326032000-ABOM-L3C_GHRSST-SSTskin-AVHRR11_D-1d_day-v02.0-fv02.0.nc,l3_file=19920326032000-ABOM-L3C_GHRSST-SSTskin-AVHRR11_D-1d_day-v02.0-fv02.0.nc,l3_source=AVHRR11_D-ABOM-L3C-v02.0,global_source=wind_source=ECMWF_interim_reanalysis,analysis_source=NCDC-L4LRblend-GLOB-AVHRR_OI,adi_source=unknown,ice_source=SSMI-NCEP-Analysis-ICE-1deg,l3_source=AVHRR11_D-ABOM-L3C-v02.0,landmask_file=lsmask.dist5.5.nc,landmask_reference=Naval Oceanographic Office (NAVOCEANO),landmask_URL=https://www.ghrsst.org/data/ghrsst-data-tools/navo-ghrsst-pp-land-sea-mask/,landmask_source=NAVOCEANO 1km Version 5.5,ice_reference=US National Weather Service - NCEP,ice_URL=http://polar.ncep.noaa.gov/seaice/Analyses.html,ice_file=19920325.ice_data.1deg.nc,ice_jdate=2448707,merge_tool=mergeL3U,mergeL3U_version=3937:3938M,quality=archive,mergeL3U_quality=archive" ;
		:references = "http://imos.org.au/sstproducts.html" ;
		:creator_url = "http://imos.org.au" ;
		:product_version = "2.0" ;
		:comment = "HRPT AVHRR experimental L3 retrieval produced by the Australian Bureau of Meteorology as a contribution to the Integrated Marine Observing System. SSTs were calibrated to drifting buoy depths (~20-30cm) followed by a cool skin correction of -0.17K to convert to a skin (~10 micron) SST. SSTs are a weighted average of the SSTs of contributing pixels (weighted by sses_standard_deviation^-2).\nWARNING: some applications are unable to properly handle signed byte values.  If byte values >127 are encountered, subtract 256 from this reported value. GRID:CONTINENTAL, SYSCODE:PRODUCTION" ;
		:Conventions = "CF-1.6" ;
		string :acknowledgment = "Any use of these data requires the following acknowledgment: \"HRPT AVHRR SSTskin retrievals were produced by the Australian Bureau of Meteorology as a contribution to the Integrated Marine Observing System - an initiative of the Australian Government being conducted as part of the National Collaborative Research Infrastructure Strategy and the Super Science Initiative.\" The imagery data were acquired from NOAA spacecraft by the Bureau, Australian Institute of Marine Science, Australian Commonwealth Scientific and Industrial Research Organization, Geoscience Australia, and Western Australian Satellite Technology and Applications Consortium." ;
		:NCO = "\"4.5.4\"" ;
data:

 lat = 19.39, 19.37, 19.35, 19.33, 19.31, 19.29, 19.27, 19.25, 19.23, 19.21, 
    19.19 ;

 lon = 70.51, 70.53, 70.55, 70.57, 70.59, 70.61, 70.63, 70.65, 70.67, 70.69, 
    70.71, 70.73, 70.75, 70.77, 70.79, 70.81, 70.83, 70.85, 70.87, 70.89, 
    70.91, 70.93, 70.95, 70.97, 70.99, 71.01 ;

 time = 354424800 ;
}

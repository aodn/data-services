netcdf imos_data_var {
dimensions:
	POSITION = 5 ;
	RANDOM = 3 ;
variables:
	double TIME ;
	double LATITUDE(POSITION) ;
	double LONGITUDE(POSITION) ;
        double DEPTH(POSITION) ;
                DEPTH:standard_name = "depth" ;
	double data_variable(POSITION) ;
		data_variable:coordinates = "TIME LATITUDE LONGITUDE DEPTH CCCC" ;
		data_variable:standard_name = "data_variable" ;
	double random_data(RANDOM) ;

// global attributes:
                :featureType = "timeSeries" ;

data:

 TIME = _ ;

 LATITUDE = _, _, _, _, _ ;

 LONGITUDE = _, _, _, _, _ ;

 DEPTH = 1, 2, 3, 4, 5 ;

 data_variable = _, _, _, _, _ ;

 random_data = _, _, _ ;
}

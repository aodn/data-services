netcdf imos_test_variable {
dimensions:
	TIME = 5 ;
	LATITUDE = 5 ;
	LONGITUDE = 5 ;
variables:
	double TIME(TIME) ;
		TIME:ancillary_variables = "TIME_quality_control" ;
	double TIME_quality_control(TIME) ;
		TIME_quality_control:standard_name = "data_variable status_flag" ;
		TIME_quality_control:quality_control_set = 1 ;
		TIME_quality_control:quality_control_conventions = "IMOS standard set using the IODE flags" ;
	double LATITUDE(LATITUDE) ;
	double LATITUDE_quality_control(TIME) ;
		LATITUDE_quality_control:standard_name = "latitude_quality_control" ;
		LATITUDE_quality_control:quality_control_set = "4" ;
		LATITUDE_quality_control:quality_control_conventions = "WOCE quality control procedure (Multidisciplinary Underway Network – CO2 measurements)" ;
	double LONGITUDE(LONGITUDE) ;
		LONGITUDE:ancillary_variables = "LONGITUDE_quality_control" ;
	double LONGITUDE_quality_control(LONGITUDE) ;
		LONGITUDE_quality_control:quality_control_set = 3 ;
		LONGITUDE_quality_control:quality_control_conventions = "very unconventional" ;
	double data_variable(TIME) ;
		data_variable:ancillary_variables = "TIME_quality_control data_variable_standard_deviation" ;
		data_variable:standard_name = "data_variable" ;
	double data_variable_standard_deviation(TIME) ;
	double data_variable1(LATITUDE) ;
		data_variable1:ancillary_variables = "LATITUDE_quality_control" ;
		data_variable1:standard_name = "data_variable1" ;
	byte bad1_quality_control ;
		bad1_quality_control:quality_control_set = 5 ;
	byte bad2_qc ;
		bad2_qc:standard_name = "data_variable status_flag" ;
	byte bad3_qc ;
		bad3_qc:quality_control_conventions = "unconventional" ;
data:

 TIME = _, _, _, _, _ ;

 TIME_quality_control = _, _, _, _, _ ;

 LATITUDE = _, _, _, _, _ ;

 LATITUDE_quality_control = _, _, _, _, _ ;

 LONGITUDE = _, _, _, _, _ ;

 LONGITUDE_quality_control = _, _, _, _, _ ;

 data_variable = _, _, _, _, _ ;

 data_variable_standard_deviation = _, _, _, _, _ ;

 data_variable1 = _, _, _, _, _ ;

 bad1_quality_control = -127 ;

 bad2_qc = -127 ;

 bad3_qc = -127 ;
}
